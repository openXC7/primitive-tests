module gtp_channel (
    input  wire          clk,
    input  wire 		 refclk_p,
    input  wire 		 refclk_n,
    input  wire          pcie_rx_n,
    input  wire          pcie_rx_p,
    output wire          pcie_tx_n,
    output wire          pcie_tx_p,
    output wire          user_led0,
    output wire          user_led1
);

wire gtrefclk0;
IBUFDS_GTE2 refclk_buffer (
	.CEB(1'd0),
	.I (refclk_p),
	.IB(refclk_n),
	.O(gtrefclk0)
);

wire gpll_lock;
wire gpll_clk;
wire gpll_refclk;
wire refclk_monitor;

(* keep *)
GTPE2_COMMON #(
	.PLL0_FBDIV(3'd5),
	.PLL0_FBDIV_45(3'd4),
	.PLL0_REFCLK_DIV(1'd1),
	.PLL1_FBDIV(3'd1),
	.PLL1_FBDIV_45(3'd5),
	.PLL1_REFCLK_DIV(2'd2)
) gtp_pll (
	.BGBYPASSB(1'd1),
	.BGPDB(1'd1),
	.BGRCALOVRD(5'd31),
	.GTREFCLK0(gtrefclk0),
	.REFCLKOUTMONITOR1(refclk_monitor),
	.PLL0LOCKEN(1'd1),
	.PLL0PD(1'd0),
	.PLL0REFCLKSEL(1'd1),
	.PLL1PD(1'd1),
	.RCALENB(1'd1),
	.PLL0LOCK      (gpll_lock),
	.PLL0OUTCLK    (gpll_clk),
	.PLL0OUTREFCLK (gpll_refclk)
);

reg  [2:0]  gtp_loopback = 3'd0;
wire        gtp_rx_init_gtrxreset0, gtp_tx_init_gttxreset0;
wire        gtp_rxphaligndone;
wire        tx_clk;
wire        rx_clk;
wire        gtp_txoutclk;
wire        gtp_rxoutclk;
reg  [19:0] gtp_txdata = 20'd0;
wire [19:0] gtp_rxdata;
reg         gtp_tx_init_txuserrdy0 = 1'd0;
reg         gtp_tx_init_txuserrdy1 = 1'd0;

reg [24:0] counter;
always @(posedge refclk_monitor) begin
	counter <= counter + 1;
end

assign user_led0 = counter[24];

GTPE2_CHANNEL #(
	// Parameters.
	.ACJTAG_DEBUG_MODE          (1'd0),
	.ACJTAG_MODE                (1'd0),
	.ACJTAG_RESET               (1'd0),
	.ADAPT_CFG0                 (1'd0),
	.ALIGN_COMMA_DOUBLE         ("FALSE"),
	.ALIGN_COMMA_ENABLE         (10'd1023),
	.ALIGN_COMMA_WORD           (2'd2),
	.ALIGN_MCOMMA_DET           ("TRUE"),
	.ALIGN_MCOMMA_VALUE         (10'd643),
	.ALIGN_PCOMMA_DET           ("TRUE"),
	.ALIGN_PCOMMA_VALUE         (9'd380),
	.CBCC_DATA_SOURCE_SEL       ("DECODED"),
	.CFOK_CFG                   (43'd5016522067584),
	.CFOK_CFG2                  (6'd32),
	.CFOK_CFG3                  (6'd32),
	.CFOK_CFG4                  (1'd0),
	.CFOK_CFG5                  (1'd0),
	.CFOK_CFG6                  (1'd0),
	.CHAN_BOND_KEEP_ALIGN       ("FALSE"),
	.CHAN_BOND_MAX_SKEW         (1'd1),
	.CHAN_BOND_SEQ_1_1          (1'd0),
	.CHAN_BOND_SEQ_1_2          (1'd0),
	.CHAN_BOND_SEQ_1_3          (1'd0),
	.CHAN_BOND_SEQ_1_4          (1'd0),
	.CHAN_BOND_SEQ_1_ENABLE     (4'd15),
	.CHAN_BOND_SEQ_2_1          (1'd0),
	.CHAN_BOND_SEQ_2_2          (1'd0),
	.CHAN_BOND_SEQ_2_3          (1'd0),
	.CHAN_BOND_SEQ_2_4          (1'd0),
	.CHAN_BOND_SEQ_2_ENABLE     (4'd15),
	.CHAN_BOND_SEQ_2_USE        ("FALSE"),
	.CHAN_BOND_SEQ_LEN          (1'd1),
	.CLK_COMMON_SWING           (1'd0),
	.CLK_CORRECT_USE            ("FALSE"),
	.CLK_COR_KEEP_IDLE          ("FALSE"),
	.CLK_COR_MAX_LAT            (4'd10),
	.CLK_COR_MIN_LAT            (4'd8),
	.CLK_COR_PRECEDENCE         ("TRUE"),
	.CLK_COR_REPEAT_WAIT        (1'd0),
	.CLK_COR_SEQ_1_1            (9'd256),
	.CLK_COR_SEQ_1_2            (1'd0),
	.CLK_COR_SEQ_1_3            (1'd0),
	.CLK_COR_SEQ_1_4            (1'd0),
	.CLK_COR_SEQ_1_ENABLE       (4'd15),
	.CLK_COR_SEQ_2_1            (9'd256),
	.CLK_COR_SEQ_2_2            (1'd0),
	.CLK_COR_SEQ_2_3            (1'd0),
	.CLK_COR_SEQ_2_4            (1'd0),
	.CLK_COR_SEQ_2_ENABLE       (4'd15),
	.CLK_COR_SEQ_2_USE          ("FALSE"),
	.CLK_COR_SEQ_LEN            (1'd1),
	.DEC_MCOMMA_DETECT          ("TRUE"),
	.DEC_PCOMMA_DETECT          ("TRUE"),
	.DEC_VALID_COMMA_ONLY       ("TRUE"),
	.DMONITOR_CFG               (12'd2560),
	.ES_CLK_PHASE_SEL           (1'd0),
	.ES_CONTROL                 (1'd0),
	.ES_ERRDET_EN               ("FALSE"),
	.ES_EYE_SCAN_EN             ("TRUE"),
	.ES_HORZ_OFFSET             (1'd0),
	.ES_PMA_CFG                 (1'd0),
	.ES_PRESCALE                (1'd0),
	.ES_QUALIFIER               (1'd0),
	.ES_QUAL_MASK               (1'd0),
	.ES_SDATA_MASK              (1'd0),
	.ES_VERT_OFFSET             (1'd0),
	.FTS_DESKEW_SEQ_ENABLE      (4'd15),
	.FTS_LANE_DESKEW_CFG        (4'd15),
	.FTS_LANE_DESKEW_EN         ("FALSE"),
	.GEARBOX_MODE               (1'd0),
	.LOOPBACK_CFG               (1'd0),
	.OUTREFCLK_SEL_INV          (2'd3),
	.PCS_PCIE_EN                ("FALSE"),
	.PCS_RSVD_ATTR              (1'd0),
	.PD_TRANS_TIME_FROM_P2      (6'd60),
	.PD_TRANS_TIME_NONE_P2      (6'd60),
	.PD_TRANS_TIME_TO_P2        (7'd100),
	.PMA_LOOPBACK_CFG           (1'd0),
	.PMA_RSV                    (10'd819),
	.PMA_RSV2                   (14'd8256),
	.PMA_RSV3                   (1'd0),
	.PMA_RSV4                   (1'd0),
	.PMA_RSV5                   (1'd0),
	.PMA_RSV6                   (1'd0),
	.PMA_RSV7                   (1'd0),
	.RXBUFRESET_TIME            (1'd1),
	.RXBUF_ADDR_MODE            ("FAST"),
	.RXBUF_EIDLE_HI_CNT         (4'd8),
	.RXBUF_EIDLE_LO_CNT         (1'd0),
	.RXBUF_EN                   ("FALSE"),
	.RXBUF_RESET_ON_CB_CHANGE   ("TRUE"),
	.RXBUF_RESET_ON_COMMAALIGN  ("FALSE"),
	.RXBUF_RESET_ON_EIDLE       ("FALSE"),
	.RXBUF_RESET_ON_RATE_CHANGE ("TRUE"),
	.RXBUF_THRESH_OVFLW         (6'd61),
	.RXBUF_THRESH_OVRD          ("FALSE"),
	.RXBUF_THRESH_UNDFLW        (3'd4),
	.RXCDRFREQRESET_TIME        (1'd1),
	.RXCDRPHRESET_TIME          (1'd1),
	.RXCDR_CFG                  (65'd19022651084486479888),
	.RXCDR_FR_RESET_ON_EIDLE    (1'd0),
	.RXCDR_HOLD_DURING_EIDLE    (1'd0),
	.RXCDR_LOCK_CFG             (4'd9),
	.RXCDR_PH_RESET_ON_EIDLE    (1'd0),
	.RXDLY_CFG                  (5'd31),
	.RXDLY_LCFG                 (6'd48),
	.RXDLY_TAP_CFG              (1'd0),
	.RXGEARBOX_EN               ("FALSE"),
	.RXISCANRESET_TIME          (1'd1),
	.RXLPMRESET_TIME            (4'd15),
	.RXLPM_BIAS_STARTUP_DISABLE (1'd0),
	.RXLPM_CFG                  (3'd6),
	.RXLPM_CFG1                 (1'd0),
	.RXLPM_CM_CFG               (1'd0),
	.RXLPM_GC_CFG               (9'd482),
	.RXLPM_GC_CFG2              (1'd1),
	.RXLPM_HF_CFG               (10'd1008),
	.RXLPM_HF_CFG2              (4'd10),
	.RXLPM_HF_CFG3              (1'd0),
	.RXLPM_HOLD_DURING_EIDLE    (1'd0),
	.RXLPM_INCM_CFG             (1'd0),
	.RXLPM_IPCM_CFG             (1'd1),
	.RXLPM_LF_CFG               (10'd1008),
	.RXLPM_LF_CFG2              (4'd10),
	.RXLPM_OSINT_CFG            (3'd4),
	.RXOOB_CFG                  (3'd6),
	.RXOOB_CLK_CFG              ("PMA"),
	.RXOSCALRESET_TIME          (2'd3),
	.RXOSCALRESET_TIMEOUT       (1'd0),
	.RXOUT_DIV                  (4'd8),
	.RXPCSRESET_TIME            (1'd1),
	.RXPHDLY_CFG                (20'd540704),
	.RXPH_CFG                   (24'd12582914),
	.RXPH_MONITOR_SEL           (1'd0),
	.RXPI_CFG0                  (1'd0),
	.RXPI_CFG1                  (1'd1),
	.RXPI_CFG2                  (1'd1),
	.RXPMARESET_TIME            (2'd3),
	.RXPRBS_ERR_LOOPBACK        (1'd0),
	.RXSLIDE_AUTO_WAIT          (3'd7),
	.RXSLIDE_MODE               ("PCS"),
	.RXSYNC_MULTILANE           (1'd0),
	.RXSYNC_OVRD                (1'd0),
	.RXSYNC_SKIP_DA             (1'd0),
	.RX_BIAS_CFG                (12'd3891),
	.RX_BUFFER_CFG              (1'd0),
	.RX_CLK25_DIV               (3'd5),
	.RX_CLKMUX_EN               (1'd1),
	.RX_CM_SEL                  (1'd1),
	.RX_CM_TRIM                 (1'd0),
	.RX_DATA_WIDTH              (5'd20),
	.RX_DDI_SEL                 (1'd0),
	.RX_DEBUG_CFG               (1'd0),
	.RX_DEFER_RESET_BUF_EN      ("TRUE"),
	.RX_DISPERR_SEQ_MATCH       ("TRUE"),
	.RX_OS_CFG                  (8'd128),
	.RX_SIG_VALID_DLY           (4'd10),
	.RX_XCLK_SEL                ("RXUSR"),
	.SAS_MAX_COM                (7'd64),
	.SAS_MIN_COM                (6'd36),
	.SATA_BURST_SEQ_LEN         (3'd5),
	.SATA_BURST_VAL             (3'd4),
	.SATA_EIDLE_VAL             (3'd4),
	.SATA_MAX_BURST             (4'd8),
	.SATA_MAX_INIT              (5'd21),
	.SATA_MAX_WAKE              (3'd7),
	.SATA_MIN_BURST             (3'd4),
	.SATA_MIN_INIT              (4'd12),
	.SATA_MIN_WAKE              (3'd4),
	.SATA_PLL_CFG               ("VCO_3000MHZ"),
	.SHOW_REALIGN_COMMA         ("TRUE"),
	.SIM_RECEIVER_DETECT_PASS   ("TRUE"),
	.SIM_RESET_SPEEDUP          ("FALSE"),
	.SIM_TX_EIDLE_DRIVE_LEVEL   ("X"),
	.SIM_VERSION                ("2.0"),
	.TERM_RCAL_CFG              (15'd16912),
	.TERM_RCAL_OVRD             (1'd0),
	.TRANS_TIME_RATE            (4'd14),
	.TST_RSV                    (1'd0),
	.TXBUF_EN                   ("TRUE"),
	.TXBUF_RESET_ON_RATE_CHANGE ("TRUE"),
	.TXDLY_CFG                  (5'd31),
	.TXDLY_LCFG                 (6'd48),
	.TXDLY_TAP_CFG              (1'd0),
	.TXGEARBOX_EN               ("FALSE"),
	.TXOOB_CFG                  (1'd0),
	.TXOUT_DIV                  (4'd8),
	.TXPCSRESET_TIME            (1'd1),
	.TXPHDLY_CFG                (20'd540704),
	.TXPH_CFG                   (11'd1920),
	.TXPH_MONITOR_SEL           (1'd0),
	.TXPI_CFG0                  (1'd0),
	.TXPI_CFG1                  (1'd0),
	.TXPI_CFG2                  (1'd0),
	.TXPI_CFG3                  (1'd0),
	.TXPI_CFG4                  (1'd0),
	.TXPI_CFG5                  (1'd0),
	.TXPI_GREY_SEL              (1'd0),
	.TXPI_INVSTROBE_SEL         (1'd0),
	.TXPI_PPMCLK_SEL            ("TXUSRCLK2"),
	.TXPI_PPM_CFG               (1'd0),
	.TXPI_SYNFREQ_PPM           (1'd1),
	.TXPMARESET_TIME            (1'd1),
	.TXSYNC_MULTILANE           (1'd0),
	.TXSYNC_OVRD                (1'd1),
	.TXSYNC_SKIP_DA             (1'd0),
	.TX_CLK25_DIV               (3'd5),
	.TX_CLKMUX_EN               (1'd1),
	.TX_DATA_WIDTH              (5'd20),
	.TX_DEEMPH0                 (1'd0),
	.TX_DEEMPH1                 (1'd0),
	.TX_DRIVE_MODE              ("DIRECT"),
	.TX_EIDLE_ASSERT_DELAY      (3'd6),
	.TX_EIDLE_DEASSERT_DELAY    (3'd4),
	.TX_LOOPBACK_DRIVE_HIZ      ("FALSE"),
	.TX_MAINCURSOR_SEL          (1'd0),
	.TX_MARGIN_FULL_0           (7'd78),
	.TX_MARGIN_FULL_1           (7'd73),
	.TX_MARGIN_FULL_2           (7'd69),
	.TX_MARGIN_FULL_3           (7'd66),
	.TX_MARGIN_FULL_4           (7'd64),
	.TX_MARGIN_LOW_0            (7'd70),
	.TX_MARGIN_LOW_1            (7'd68),
	.TX_MARGIN_LOW_2            (7'd66),
	.TX_MARGIN_LOW_3            (7'd64),
	.TX_MARGIN_LOW_4            (7'd64),
	.TX_PREDRIVER_MODE          (1'd0),
	.TX_RXDETECT_CFG            (13'd6194),
	.TX_RXDETECT_REF            (3'd4),
	.TX_XCLK_SEL                ("TXOUT"),
	.UCODEER_CLR                (1'd0),
	.USE_PCS_CLK_PHASE_SEL      (1'd0)
) GTPE2_CHANNEL (
	// Inputs.
	.CFGRESET             (1'd0),
	.CLKRSVD0             (1'd0),
	.CLKRSVD1             (1'd0),
	.DMONFIFORESET        (1'd0),
	.DMONITORCLK          (1'd0),
	.DRPADDR              (),
	.DRPCLK               (),
	.DRPDI                (),
	.DRPEN                (1'b0),
	.DRPWE                (),
	.EYESCANMODE          (1'd0),
	.EYESCANRESET         (1'd0),
	.EYESCANTRIGGER       (1'd0),
	.GTPRXN               (pcie_rx_n),
	.GTPRXP               (pcie_rx_p),
	.GTRESETSEL           (1'd0),
	.GTRSVD               (1'd0),
	.GTRXRESET            (gtp_rx_init_gtrxreset0),
	.GTTXRESET            (gtp_tx_init_gttxreset0),
	.LOOPBACK             (gtp_loopback),
	.PCSRSVDIN            (1'd0),
	.PLL0CLK              (gpll_clk),
	.PLL0REFCLK           (gpll_refclk),
	.PLL1CLK              (1'd0),
	.PLL1REFCLK           (1'd0),
	.PMARSVDIN0           (1'd0),
	.PMARSVDIN1           (1'd0),
	.PMARSVDIN2           (1'd0),
	.PMARSVDIN3           (1'd0),
	.PMARSVDIN4           (1'd0),
	.RESETOVRD            (1'd0),
	.RX8B10BEN            (1'd0),
	.RXADAPTSELTEST       (1'd0),
	.RXBUFRESET           (1'd0),
	.RXCDRFREQRESET       (1'd0),
	.RXCDRHOLD            (1'd0),
	.RXCDROVRDEN          (1'd0),
	.RXCDRRESET           (1'd0),
	.RXCDRRESETRSV        (1'd0),
	.RXCHBONDEN           (1'd0),
	.RXCHBONDI            (1'd0),
	.RXCHBONDLEVEL        (1'd0),
	.RXCHBONDMASTER       (1'd0),
	.RXCHBONDSLAVE        (1'd0),
	.RXCOMMADETEN         (1'd1),
	.RXDDIEN              (1'd1),
	.RXDFEXYDEN           (1'd0),
	.RXDLYBYPASS          (1'd0),
	.RXDLYEN              (1'd0),
	.RXDLYOVRDEN          (1'd0),
	.RXDLYSRESET          (1'b0),
	.RXELECIDLEMODE       (2'd3),
	.RXGEARBOXSLIP        (1'd0),
	.RXLPMHFHOLD          (1'd0),
	.RXLPMHFOVRDEN        (1'd0),
	.RXLPMLFHOLD          (1'd0),
	.RXLPMLFOVRDEN        (1'd0),
	.RXLPMOSINTNTRLEN     (1'd0),
	.RXLPMRESET           (1'd0),
	.RXMCOMMAALIGNEN      (1'd0),
	.RXOOBRESET           (1'd0),
	.RXOSCALRESET         (1'd0),
	.RXOSHOLD             (1'd0),
	.RXOSINTCFG           (2'd2),
	.RXOSINTEN            (1'd1),
	.RXOSINTHOLD          (1'd0),
	.RXOSINTID0           (1'd0),
	.RXOSINTNTRLEN        (1'd0),
	.RXOSINTOVRDEN        (1'd0),
	.RXOSINTPD            (1'd0),
	.RXOSINTSTROBE        (1'd0),
	.RXOSINTTESTOVRDEN    (1'd0),
	.RXOSOVRDEN           (1'd0),
	.RXOUTCLKSEL          (2'd2),
	.RXPCOMMAALIGNEN      (1'd0),
	.RXPCSRESET           (1'd0),
	.RXPD                 (2'b00),
	.RXPHALIGN            (1'd0),
	.RXPHALIGNEN          (1'd0),
	.RXPHDLYPD            (1'd0),
	.RXPHDLYRESET         (1'd0),
	.RXPHOVRDEN           (1'd0),
	.RXPMARESET           (1'd0),
	.RXPOLARITY           (1'd0),
	.RXPRBSCNTRESET       (1'd0),
	.RXPRBSSEL            (1'd0),
	.RXRATE               (1'd0),
	.RXRATEMODE           (1'd0),
	.RXSLIDE              (1'd0),
	.RXSYNCALLIN          (gtp_rxphaligndone),
	.RXSYNCIN             (1'd0),
	.RXSYNCMODE           (1'd1),
	.RXSYSCLKSEL          (1'd0),
	.RXUSERRDY            (1'b1),
	.RXUSRCLK             (rx_clk),
	.RXUSRCLK2            (rx_clk),
	.SETERRSTATUS         (1'd0),
	.SIGVALIDCLK          (1'd0),
	.TSTIN                (20'd1048575),
	.TX8B10BBYPASS        (1'd0),
	.TX8B10BEN            (1'd0),
	.TXBUFDIFFCTRL        (3'd4),
	.TXCHARDISPMODE       ({gtp_txdata[19], gtp_txdata[9]}),
	.TXCHARDISPVAL        ({gtp_txdata[18], gtp_txdata[8]}),
	.TXCHARISK            (1'd0),
	.TXCOMINIT            (1'd0),
	.TXCOMSAS             (1'd0),
	.TXCOMWAKE            (1'd0),
	.TXDATA               ({gtp_txdata[17:10], gtp_txdata[7:0]}),
	.TXDEEMPH             (1'd0),
	.TXDETECTRX           (1'd0),
	.TXDIFFCTRL           (4'd8),
	.TXDIFFPD             (1'd0),
	.TXDLYBYPASS          (1'd1),
	.TXDLYEN              (1'd0),
	.TXDLYHOLD            (1'd0),
	.TXDLYOVRDEN          (1'd0),
	.TXDLYSRESET          (1'b0),
	.TXDLYUPDOWN          (1'd0),
	.TXELECIDLE           (1'd0),
	.TXHEADER             (1'd0),
	.TXINHIBIT            (1'b0),
	.TXMAINCURSOR         (1'd0),
	.TXMARGIN             (1'd0),
	.TXOUTCLKSEL          (2'd2),
	.TXPCSRESET           (1'd0),
	.TXPD                 (1'd0),
	.TXPDELECIDLEMODE     (1'd0),
	.TXPHALIGN            (1'b0),
	.TXPHALIGNEN          (1'd0),
	.TXPHDLYPD            (1'd0),
	.TXPHDLYRESET         (1'd0),
	.TXPHDLYTSTCLK        (1'd0),
	.TXPHINIT             (1'b0),
	.TXPHOVRDEN           (1'd0),
	.TXPIPPMEN            (1'd0),
	.TXPIPPMOVRDEN        (1'd0),
	.TXPIPPMPD            (1'd0),
	.TXPIPPMSEL           (1'd1),
	.TXPIPPMSTEPSIZE      (1'd0),
	.TXPISOPD             (1'd0),
	.TXPMARESET           (1'd0),
	.TXPOLARITY           (1'd0),
	.TXPOSTCURSOR         (1'd0),
	.TXPOSTCURSORINV      (1'd0),
	.TXPRBSFORCEERR       (1'd0),
	.TXPRBSSEL            (1'd0),
	.TXPRECURSOR          (1'd0),
	.TXPRECURSORINV       (1'd0),
	.TXRATE               (1'd0),
	.TXRATEMODE           (1'd0),
	.TXSEQUENCE           (1'd0),
	.TXSTARTSEQ           (1'd0),
	.TXSWING              (1'd0),
	.TXSYNCALLIN          (1'd0),
	.TXSYNCIN             (1'd0),
	.TXSYNCMODE           (1'd0),
	.TXSYSCLKSEL          (1'd0),
	.TXUSERRDY            (gtp_tx_init_txuserrdy0),
	.TXUSRCLK             (tx_clk),
	.TXUSRCLK2            (tx_clk),

	// Outputs.
	.DMONITOROUT          (),
	.DRPDO                (),
	.DRPRDY               (),
	.EYESCANDATAERROR     (),
	.GTPTXN               (pcie_tx_n),
	.GTPTXP               (pcie_tx_p),
	.PCSRSVDOUT           (),
	.PHYSTATUS            (),
	.PMARSVDOUT0          (),
	.PMARSVDOUT1          (),
	.RXBUFSTATUS          (),
	.RXBYTEISALIGNED      (),
	.RXBYTEREALIGN        (),
	.RXCDRLOCK            (),
	.RXCHANBONDSEQ        (),
	.RXCHANISALIGNED      (),
	.RXCHANREALIGN        (),
	.RXCHARISCOMMA        (),
	.RXCHARISK            ({gtp_rxdata[18], gtp_rxdata[8]}),
	.RXCHBONDO            (),
	.RXCLKCORCNT          (),
	.RXCOMINITDET         (),
	.RXCOMMADET           (),
	.RXCOMSASDET          (),
	.RXCOMWAKEDET         (),
	.RXDATA               ({gtp_rxdata[17:10], gtp_rxdata[7:0]}),
	.RXDATAVALID          (),
	.RXDISPERR            ({gtp_rxdata[19], gtp_rxdata[9]}),
	.RXDLYSRESETDONE      (),
	.RXELECIDLE           (),
	.RXHEADER             (),
	.RXHEADERVALID        (),
	.RXNOTINTABLE         (),
	.RXOSINTDONE          (),
	.RXOSINTSTARTED       (),
	.RXOSINTSTROBEDONE    (),
	.RXOSINTSTROBESTARTED (),
	.RXOUTCLK             (gtp_rxoutclk),
	.RXOUTCLKFABRIC       (),
	.RXOUTCLKPCS          (),
	.RXPHALIGNDONE        (gtp_rxphaligndone),
	.RXPHMONITOR          (),
	.RXPHSLIPMONITOR      (),
	.RXPMARESETDONE       (),
	.RXPRBSERR            (),
	.RXRATEDONE           (),
	.RXRESETDONE          (),
	.RXSTARTOFSEQ         (),
	.RXSTATUS             (),
	.RXSYNCDONE           (),
	.RXSYNCOUT            (),
	.RXVALID              (),
	.TXBUFSTATUS          (),
	.TXCOMFINISH          (),
	.TXDLYSRESETDONE      (),
	.TXGEARBOXREADY       (),
	.TXOUTCLK             (gtp_txoutclk),
	.TXOUTCLKFABRIC       (),
	.TXOUTCLKPCS          (),
	.TXPHALIGNDONE        (),
	.TXPHINITDONE         (),
	.TXPMARESETDONE       (),
	.TXRATEDONE           (),
	.TXRESETDONE          (),
	.TXSYNCDONE           (),
	.TXSYNCOUT            ()
);


endmodule
